--Bibliotecas
library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity NAND2Gate is
	port( input0 : in std_logic;
			input1 : in std_logic;
			output : out std_logic
	);
end NAND2Gate;

architecture Structural of NAND2Gate is

	signal s_andOut : std_logic;

begin 

	and_gate : entity work.AND2Gate(Behavioral)
							port map (  input0 => input0,
											input1 => input1,
											output => s_andOut);
	
	not_gate : entity work.NOTGate(Behavioral)
							port map (  input => s_andOut,
											output => output);
end Structural;